//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//
// Description: 
//
//----------------------------------------------------------------------
//
// Device:
// Block:       
// Designer:    Martin Marinov
//
//----------------------------------------------------------------------
//
// $URL:$
// $Revision:$
// $Date:$
// $Author:$
//
//----------------------------------------------------------------------
`default_nettype none

module sync_reg_2edge #(
    parameter                               SYNC_REG_WDTH   = 1
) (
                            input wire                              clk1,
                            input wire                              clk2,
                            input wire [SYNC_REG_WDTH-1         :0] sync_sig,
(* ASYNC_REG = "TRUE" *)    output reg [SYNC_REG_WDTH-1         :0] sync_reg1
);

//*****************************************************************************
// Local defines
//*****************************************************************************
(* ASYNC_REG = "TRUE" *)    reg [SYNC_REG_WDTH-1      :0] sync_reg0 = {SYNC_REG_WDTH{1'b0}};
//(* ASYNC_REG = "TRUE" *)    reg [SYNC_REG_WDTH-1      :0] sync_reg1;

//*****************************************************************************
// CDC sync
//*****************************************************************************


    always @(posedge clk1) begin
        sync_reg0 <= sync_sig;
    end

    always @(posedge clk2) begin
        sync_reg1 <= sync_reg0;
    end


//*****************************************************************************
// Output assignments
//*****************************************************************************
//assign synced_sig = sync_reg1;


//*****************************************************************************
//                                  END OF FILE
//*****************************************************************************
endmodule

`resetall
